* C:\Users\mistr\eSim-Workspace\decoder\decoder.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/14/21 21:59:07

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U6  Net-_U3-Pad3_ Net-_U3-Pad4_ Net-_U10-Pad1_ d_and		
U7  Net-_U3-Pad3_ Net-_U4-Pad2_ Net-_U10-Pad2_ d_and		
U9  Net-_U5-Pad2_ Net-_U3-Pad4_ Net-_U10-Pad3_ d_and		
U8  Net-_U5-Pad2_ Net-_U4-Pad2_ Net-_U10-Pad4_ d_and		
U10  Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad3_ Net-_U10-Pad4_ Y3 Y2 Y1 Y0 dac_bridge_4		
R1  Y3 ? 100		
R4  Y2 GND 100		
R2  Y1 GND 100		
U3  A1 A0 Net-_U3-Pad3_ Net-_U3-Pad4_ adc_bridge_2		
v1  A1 GND DC		
v2  A0 GND DC		
U1  A1 plot_v1		
U2  A0 plot_v1		
U4  Net-_U3-Pad4_ Net-_U4-Pad2_ d_inverter		
U5  Net-_U3-Pad3_ Net-_U5-Pad2_ d_inverter		
R3  Y0 GND 100		
U12  Y3 plot_v1		
U14  Y2 plot_v1		
U11  Y0 plot_v1		
U13  Y1 plot_v1		

.end
